module invert ( 
    input wire i, 
    output wire o 
); 

assign o = !i; 
endmodule 

module and2 ( 
    input wire i0, i1, 
    output wire o 
); 

assign o = i0 & i1; 
endmodule 

module or2 ( 
    input wire i0, i1, 
    output wire o
); 

assign o = i0 | i1; 
endmodule 

module xor2 ( 
    input wire i0, i1, 
    output wire o 
); 

assign o = i0 ^ i1; 
endmodule 

module nand2 ( 
    input wire i0, i1, 
    output wire o 
); 
    
wire t;

and2 and2_0 ( i0, i1, t); 
invert invert_0 ( t, o); 
endmodule 

module nor2 ( 
    input wire i0, i1, 
    output wire o 
); 

wire t; or2 or2_0 ( i0, i1, t); 
invert invert_0 ( t, o ); 
endmodule 

module xnor2 ( 
    input wire i0, i1, 
    output wire o 
); 

wire t; 
xor2 xor2_0 ( i0, i1, t ); 
invert invert_0 ( t, o ); 
endmodule 

module and3 ( 
    input wire i0, i1, i2, 
    output wire o 
); 

wire t; and2 and2_0 ( i0, i1, t ); 
and2 and2_1 ( i2, t, o ); 
endmodule 

module or3 ( 
    input wire i0, i1, i2, 
    output wire o 
); 

wire t; 
or2 or2_0 ( i0, i1, t ); 
or2 or2_1 ( i2, t, o ); 
endmodule 

module nor3 ( 
    input wire i0, i1, i2, 
    output wire o 
); 
wire t; 
or2 or2_0 ( i0, i1, t ); 
nor2 nor2_0 ( i2, t, o); 
endmodule 

module nand3 ( 
    input wire i0, i1, i2, 
    output wire o 
); 
wire t; 
and2 and2_0 ( i0, i1, t ); 
nand2 nand2_1 ( i2, t, o ); 
endmodule 

module xor3 ( 
    input wire i0, i1, i2, 
    output wire o 
); 

wire t; 
xor2 xor2_0 ( i0, i1, t ); 
xor2 xor2_1 ( i2, t, o );
endmodule
 
module xnor3 ( 
    input wire i0, i1, i2, 
    output wire o 
); 

wire t; 
xor2 xor2_0 ( i0, i1, t ); 
xnor2 xnor2_0 ( i2, t, o ); 
endmodule 

module mux2 ( 
    input wire i0, i1, j, 
    output wire o 
); 

assign o = (j == 0) ? i0 : i1; 
endmodule 

module mux4 ( 
    input wire [0:3] i, 
    input wire j1, j0, 
    output wire o 
); 

wire t0, t1; 
mux2 mux2_0 ( i[0], i[1], j1, t0 ); 
mux2 mux2_1 ( i[2], i[3], j1, t1 ); 
mux2 mux2_2 ( t0, t1, j0, o ); 
endmodule 

module mux8 ( 
    input wire [0:7] i, 
    input wire j2, j1, j0, 
    output wire o 
); 

wire t0, t1; 
mux4 mux4_0 ( i[0:3], j2, j1, t0 );
 mux4 mux4_1 ( i[4:7], j2, j1, t1 ); 
 mux2 mux2_0 (t0, t1, j0, o ); 
endmodule